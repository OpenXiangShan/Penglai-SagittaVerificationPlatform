`ifndef TCNT_APB_MASTER_PKG__SV
`define TCNT_APB_MASTER_PKG__SV

package tcnt_apb_master_pkg;
	import uvm_pkg::*;
    import tcnt_apb_dec::*;

	`include "tcnt_apb_master_agent_cfg.sv"
	`include "tcnt_apb_master_agent_transaction.sv"
	`include "tcnt_apb_master_agent_sequence.sv"
	`include "tcnt_apb_master_agent_sequencer.sv"
    `include "tcnt_apb_master_agent_driver_callback.sv"
	`include "tcnt_apb_master_agent_driver.sv"
	`include "tcnt_apb_master_agent_monitor.sv"
	`include "tcnt_apb_master_agent.sv"
endpackage:tcnt_apb_master_pkg
import tcnt_apb_master_pkg::*;

`endif
